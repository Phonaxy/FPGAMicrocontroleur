--Question a.1.1
--Pour calculer C en fonction de A et B on a besoin d'un AND 
--Pour calculer S en fonction de A et B on a besoin d'un XOR
	
--Question a.1.2
